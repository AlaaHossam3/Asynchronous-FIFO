package shared_pkg;

int error_count   = 0;
int correct_count = 0;
bit test_finished;
event trigger;
    
endpackage